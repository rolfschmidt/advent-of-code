module main

fn main() {
	println(day17a())
	println(day17b())
}
