module main

fn main() {
	println(day15a())
	println(day15b())
}
