module main

fn test_day03a() {
	assert day03a() == 164
}

fn test_day03b() {
	assert day03b() == 5007658656
}
