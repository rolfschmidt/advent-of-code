module main

fn test_day20a() {
	assert day20a() == 111936085519519
}

fn test_day20b() {
	assert day20b() == 1792
}
