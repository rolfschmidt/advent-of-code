module main

fn main() {
	println(day18a())
	println(day18b())
}
