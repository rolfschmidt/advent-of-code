module main

fn main() {
	println('Part 1:')
	println('Day 1: $day01a()')
	println('Day 2: $day02a()')
	println('Day 3: $day03a()')
	println('Day 4: $day04a()')
	println('Day 5: $day05a()')
	println('Day 6: $day06a()')
	println('Day 7: $day07a()')
	println('Day 8: $day08a()')
	println('Day 9: $day09a()')
	println('Day 10: $day10a()')
	println('Day 11: $day11a()')
	println('Day 12: $day12a()')
	println('Day 13: $day13a()')
	println('Day 14: $day14a()')
	println('Day 15: $day15a()')
	println('Day 16: $day16a()')
	println('Day 17: $day17a()')
	println('Day 18: $day18a()')
	println('Day 19: $day19a()')
	println('Day 20: $day20a()')
	println('Day 21: $day21a()')
	println('Day 22: $day22a()')
	println('Day 23: $day23a()')
	println('Day 24: $day24a()')
	println('Day 25: $day25a()')
	// println('Part 2:')
	// println('Day 1: ${day01b()}')
	// println('Day 2: ${day02b()}')
	// println('Day 3: ${day03b()}')
	// println('Day 4: ${day04b()}')
	// println('Day 5: ${day05b()}')
	// println('Day 6: ${day06b()}')
	// println('Day 7: ${day07b()}')
	// println('Day 8: ${day08b()}')
	// println('Day 9: ${day09b()}')
	// println('Day 10: ${day10b()}')
	// println('Day 11: ${day11b()}')
	// println('Day 12: ${day12b()}')
	// println('Day 13: ${day13b()}')
	// println('Day 14: ${day14b()}')
	// println('Day 15: ${day15b()}')
	// println('Day 16: ${day16b()}')
	// println('Day 17: ${day17b()}')
	// println('Day 18: ${day18b()}')
	// println('Day 19: ${day19b()}')
	// println('Day 20: ${day20b()}')
	// println('Day 21: ${day21b()}')
	// println('Day 22: ${day22b()}')
	// println('Day 23: ${day23b()}')
	// println('Day 24: ${day24b()}')
	// println('Day 25: ${day25b()}')
}
