module main

fn main() {
    println(day01a())
    println(day01b())

}