module main

fn test_day25a() {
	assert day25a() == 16933668
}

fn test_day25b() {
	assert day25b() == 0
}
