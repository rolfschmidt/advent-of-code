module main

fn test_day16a() {
	assert day16a() == 29759
}

fn test_day16b() {
	assert day16b() == 1307550234719
}
