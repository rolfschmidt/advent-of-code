module main

fn test_day01a() {
    assert day01a() == 858496
}

fn test_day01b() {
    assert day01b() == 263819430
}
