module main

fn test_day12a() {
	assert day12a() == 1838
}

fn test_day12b() {
	assert day12b() == 89936
}
