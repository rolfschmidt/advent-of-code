module main

fn test_day02a() {
    assert day02a() == 586
}

fn test_day02b() {
    assert day02b() == 352
}
