module main

fn test_day21a() {
	assert day21a() == '1930'
}

fn test_day21b() {
	assert day21b() == 'spcqmzfg,rpf,dzqlq,pflk,bltrbvz,xbdh,spql,bltzkxx'
}
