module main

fn main() {
	println(day10a())
	println(day10b())
}
