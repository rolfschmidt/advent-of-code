module main

fn test_day01a() {
    assert day01a() == 437931
}

fn test_day01b() {
    assert day01b() == 157667328
}
