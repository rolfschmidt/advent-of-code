module main

fn test_day10a() {
	assert day10a() == 2760
}

fn test_day10b() {
	assert day10b() == 13816758796288
}
