module main

fn test_day14a() {
	assert day14a() == 3059488894985
}

fn test_day14b() {
	assert day14b() == 0
}
