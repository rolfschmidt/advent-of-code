module main

fn test_day06a() {
	assert day06a() == 6443
}

fn test_day06b() {
	assert day06b() == 3232
}
