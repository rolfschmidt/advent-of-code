module main

fn main() {
	println(day11a())
	println(day11b())
}
