module main

fn test_day09a() {
	assert day09a() == 3199139634
}

fn test_day09b() {
	assert day09b() == 438559930
}
