module main

fn test_day22a() {
	assert day22a() == 30780
}

fn test_day22b() {
	// assert day22b() == 36621
}
