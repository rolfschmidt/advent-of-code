module main

fn main() {
	println(day23a())
	println(day23b())
}
