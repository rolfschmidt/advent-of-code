module main

fn main() {
	println(day04a())
	println(day04b())
}
