module main

fn test_day11a() {
	// assert day11a() == 2222
}

fn test_day11b() {
	// assert day11b() == 2032
}
