module main

fn test_day05a() {
	assert day05a() == 874
}

fn test_day05b() {
	assert day05b() == 594
}
