module main

fn main() {
	println(day13a())
	println(day13b())
}
