module main

fn main() {
	println(day05a())
	println(day05b())
}
