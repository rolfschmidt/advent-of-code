module main

fn main() {
	println(day20a())
	println(day20b())
}
