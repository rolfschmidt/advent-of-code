module main

fn test_day23a() {
	assert day23a() == '32658947'
}

fn test_day23b() {
	// assert day23b() == '683486010900'
}
