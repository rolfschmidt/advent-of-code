module main

fn main() {
	println(day12a())
	println(day12b())
}
