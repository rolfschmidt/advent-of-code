module main

fn main() {
	println(day22a())
	println(day22b())
}
