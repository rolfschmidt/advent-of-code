module main

fn main() {
	println(day14a())
	println(day14b())
}
