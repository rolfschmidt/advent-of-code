module main

fn test_day17a() {
	assert day17a() == 322
}

fn test_day17b() {
	// assert day17b() == 2000
}
