module main

fn main() {
	println(day08a())
	println(day08b())
}
