module main

fn test_day19a() {
	assert day19a() == 132
}

fn test_day19b() {
	assert day19b() == 306
}
