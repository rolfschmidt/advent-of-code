module main

fn main() {
	println(day25a())
	println(day25b())
}
