module main

fn test_day07a() {
	assert day07a() == 378
}

fn test_day07b() {
	assert day07b() == 27526
}
