module main

fn main() {
	println(day21a())
	println(day21b())
}
