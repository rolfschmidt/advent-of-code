module main

fn main() {
    println(day02a())
    println(day02b())
}