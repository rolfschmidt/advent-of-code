module main

fn test_day24a() {
	assert day24a() == 275
}

fn test_day24b() {
	assert day24b() == 3537
}
