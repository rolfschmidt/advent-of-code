module main

fn main() {
	println(day09a())
	println(day09b())
}
