module main

fn main() {
	println(day16a())
	println(day16b())
}
