module main

fn main() {
	println(day24a())
	println(day24b())
}
