module main

fn test_bindec() {
	assert bindec('000000000000000000000000000000001011') == 11
	assert bindec('000000000000000000000000000001001001') == 73
	assert bindec('000000000000000000000000000001000000') == 64
	assert bindec('000000000000010011100011111010011011') == 5127835
	assert bindec('000000000000100101000100010110001111') == 9717135
	assert bindec('110000001000100111101100000100001000') == 51684229384
}

fn test_decbin() {
	assert decbin(11, 36) == '000000000000000000000000000000001011'
	assert decbin(73, 36) == '000000000000000000000000000001001001'
	assert decbin(64, 36) == '000000000000000000000000000001000000'
	assert decbin(5127835, 36) == '000000000000010011100011111010011011'
	assert decbin(9717135, 36) == '000000000000100101000100010110001111'
	assert decbin(51684229384, 36) == '110000001000100111101100000100001000'
}
