module main

fn test_day08a() {
	assert day08a() == 1475
}

fn test_day08b() {
	assert day08b() == 1270
}
