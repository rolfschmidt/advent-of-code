module main

fn test_day13a() {
	assert day13a() == 410
}

fn test_day13b() {
	assert day13b() == 600691418730595
}
