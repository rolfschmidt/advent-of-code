module main

fn main() {
	println(day19a())
	println(day19b())
}
