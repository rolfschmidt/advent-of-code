module main

fn main() {
	println(day06a())
	println(day06b())
}
