module main

fn main() {
	println(day03a())
	println(day03b())
}
