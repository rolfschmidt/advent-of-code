module main

fn main() {
	println(day07a())
	println(day07b())
}
