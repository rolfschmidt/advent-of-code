module main

fn test_day04a() {
	assert day04a() == 222
}

fn test_day04b() {
	assert day04b() == 140
}
